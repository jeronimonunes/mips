module ula(inputA, inputB, operation, outputA);

input [32:0] inputA;
input [32:0] inputB;
//TODO Find number of operation bits on mips
input operation;
output reg [32:0] outputA;


endmodule
